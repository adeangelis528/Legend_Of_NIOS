module sprite_rom ( input [5:0]	addr,
						output [31:0]	data
					 );

	parameter ADDR_WIDTH = 5;
   parameter DATA_WIDTH =  32;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  //Wall Tile
        32'b11111111111111111111111111111111,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b11111111111111111111111111111111,
		  
		  //Floor Tile
		  32'b00000000000000000000000000000000,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b01111111111111111111111111111110,
		  32'b00000000000000000000000000000000,
        };

	assign data = ROM[addr];

endmodule  