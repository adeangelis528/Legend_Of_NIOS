/*
Modified sprite table ROM
takes the input of DrawX and DrawY and returns
if a floor or wall should be drawn
1 = draw wall
0 = draw floor
MAKE SURE DOORS MATCH UP
*/
module level_rom ( input [9:0]	DrawX, DrawY,
						 input logic [2:0] room,
						 output logic bg_type
					 );

	logic [19:0] data;
	
	// ROM definition		
	//Each room contains 20x15 background tiles
	parameter [0:119][19:0] ROM = {
	     //Room 0
		  20'b00000000000000000000,
		  20'b11111111100111111111,
		  20'b10000000000000000001,
        20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000000,
		  20'b10000000000000000000,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111,
		  
		  //Room 1
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10000000000000000001,
		  20'b10000000011000000001,
		  20'b10000000011000000001,
		  20'b10000000011000000001,
		  20'b00001111111111110000,
		  20'b00001111111111110000,
		  20'b10000000011000000001,
		  20'b10000000011000000001,
		  20'b10000000011000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111,
		  
		  //Room 2
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10111111000011111101,
		  20'b10100000000000000101,
		  20'b10100000000000000101,
		  20'b10100000000000000101,
		  20'b10100110000001100101,
		  20'b10100110000001100101,
		  20'b10100000000000000101,
		  20'b10100000000000000101,
		  20'b10100000000000000101,
		  20'b10111111000011111101,
		  20'b10000000000000000001,
		  20'b11111111100111111111,
		  
		  //Room 3
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10000000000000000001,
		  20'b10011111111111111001,
		  20'b10010000000000000001,
		  20'b10010000000000000001,
		  20'b00010011111111111111,
		  20'b00010000000000000001,
		  20'b11110000000000000001,
		  20'b11111111111111111001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b11111111100111111111,
		  
		  //Room 4
		  20'b00000000000000000000,
		  20'b11111111100111111111,
		  20'b10000000000000000001,
        20'b10010000000000000001,
		  20'b10111000000000000001,
		  20'b10010000000001000001,
		  20'b10000000000011100001,
		  20'b10000000000001000000,
		  20'b10000001000000000000,
		  20'b10000011100000000001,
		  20'b10000001000010000001,
		  20'b10000000000111000001,
		  20'b10000000000010000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111,
		  
		  //Room 5
		  20'b00000000000000000000,
		  20'b11111111100111111111,
		  20'b10000000000000000001,
        20'b10000000000000000001,
		  20'b10000000011000000001,
		  20'b10000000111100000001,
		  20'b10000001111110000001,
		  20'b00000011111111000000,
		  20'b00000011111111000000,
		  20'b10000001111110000001,
		  20'b10000000111100000001,
		  20'b10000000011000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111,
		  
		  //Room 6
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10110000000000001101,
		  20'b10100000000000000101,
		  20'b10000000000000000001,
		  20'b10000110000001100001,
		  20'b10000100000000100001,
		  20'b10000100000000100001,
		  20'b10000110000001100001,
		  20'b10000000000000000001,
		  20'b10100000000000000101,
		  20'b10110000000000001101,
		  20'b10000000000000000001,
		  20'b11111111100111111111,
		  
		  //Room 7
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10000001010111010101,
		  20'b10000001010101011101,
		  20'b10000001010101001001,
		  20'b10000001110111001001,
		  20'b00000000000000000001,
		  20'b00000000000000000001,
		  20'b10100101010001000001,
		  20'b10101101010001000001,
		  20'b10110101010101000001,
		  20'b10100101011011000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111
        };

	always_comb begin
		  
		data = ROM[15 * room + (DrawY/32)];
		bg_type = data[DrawX/32];
	
	end

endmodule