module sprite_rom ( input [6:0]	addr,
						output [31:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  32;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  //Wall Tile, code 0
        32'b11111111111111111111111111111111,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b11111111111111111111111111111111,
		  
		  //Floor Tile, code 1
		  32'b00000000000000000000000000000000,
		  32'b00000111111111111111111111100000,
		  32'b00011111111111111111111111111000,
		  32'b00100000000000000000000000000100,
		  32'b00101111111111111111111111110100,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b00101111111111111111111111110100,
		  32'b00100000000000000000000000000100,
		  32'b00011111111111111111111111111000,
		  32'b00000111111111111111111111100000,
		  32'b00000000000000000000000000000000,
		  
		  //Player Character, code 2
		  32'b11000000000000000000000000000011,
		  32'b10000000000000111100000000000001,
		  32'b00000000000001111110000000000000,
		  32'b00000000000000111100000000000000,
		  32'b00000000000010011001000000000000,
		  32'b00000000000001011010000000000000,
		  32'b00000000000000111100000000000000,
		  32'b00000000000000011000000000000000,
		  32'b00000000000000011000000000000000,
		  32'b00000000000000011000000000000000,
		  32'b00000000000000011000000000000000,
		  32'b00000000000000100100000000000000,
		  32'b00000000000001000010000000000000,
		  32'b00000000000010000001000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b00000000000000000000000000000000,
		  32'b10000000000000000000000000000001,
		  32'b11000000000000000000000000000011,
		  
		  //Unused
		  32'b11111111111111111111111111111111,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b11111111111111111111111111111111
        };

	assign data = ROM[addr];

endmodule  