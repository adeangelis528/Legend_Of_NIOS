//-------------------------------------------------------------------------
//      Legend of NIOS                                                   --
//      Andrew DeAngelis, Michael Recklein                               --
//      Fall 2017                                                        --
//                                                                       --
//      Built on Lab 8 USB interface                                     --
//                                                                       --
//                                                                       --
//-------------------------------------------------------------------------


module lab8( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1,
             // VGA Interface 
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK      //SDRAM Clock
                    );
    
    logic Reset_h, Clk;
    logic [15:0] keycode;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs;
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),    
                            .OTG_RST_N(OTG_RST_N)
    );
     
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     nios_system nios_system(
                             .clk_clk(Clk),         
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_out_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w),
									  .entity_active_export(toNIOS_Active),
									  .entity_dir_export(sel_dir),
									  .entity_read_export(read),
									  .entity_select_export(select),
									  .entity_write_export(write),
									  .entity_x_export(toNIOS_X),
									  .entity_y_export(toNIOS_Y),
									  .entity_type_export(toNIOS_Type)
    );
  
    // Use PLL to generate the 25MHZ VGA_CLK. Do not modify it.
    // vga_clk vga_clk_instance(
    //     .clk_clk(Clk),
    //     .reset_reset_n(1'b1),
    //     .altpll_0_c0_clk(VGA_CLK),
    //     .altpll_0_areset_conduit_export(),    
    //     .altpll_0_locked_conduit_export(),
    //     .altpll_0_phasedone_conduit_export()
    // );
	 
    always_ff @ (posedge Clk) begin
        if(Reset_h)
            VGA_CLK <= 1'b0;
        else
            VGA_CLK <= ~VGA_CLK;
    end
    
	 //Extra logic for graphical interconnections
	 logic[9:0] DrawX, DrawY;
	 logic[9:0] Player_X, Player_Y;
	 logic[7:0] bg_r, bg_g, bg_b;
	 logic[10:0] font_addr;
	 logic[3:0] text_offset;
	 logic draw_text, bg_type;
	 logic[2:0] room, doorcode;
	 logic[1:0] health;
	 logic[3:0] score1, score2;
	 
	 //Temporary
	 //assign room = 0;
	 //assign bg_type = 0;
	   logic[2:0] select;
	   logic read, write, initialize;
	   logic[2:0] sel_dir;
	   logic[9:0] Enemy1_X, Enemy2_X, Enemy3_X, Enemy4_X, Enemy5_X;
	   logic[9:0] Enemy1_Y, Enemy2_Y, Enemy3_Y, Enemy4_Y, Enemy5_Y;
	   logic Enemy1_Active, Enemy2_Active, Enemy3_Active, Enemy4_Active, Enemy5_Active;
		logic Damage_E1, Damage_E2, Damage_E3, Damage_E4, Damage_E5;
		logic[1:0] Type_E1, Type_E2, Type_E3, Type_E4, Type_E5;
	   logic[9:0] toNIOS_X, toNIOS_Y;
		logic[1:0] toNIOS_Type;
	   logic[2:0] toEnemy1_dir, toEnemy2_dir, toEnemy3_dir, toEnemy4_dir, toEnemy5_dir;
	   logic toNIOS_Active;
		logic game_over, player_attack, game_reset;
		
		assign game_reset = game_over | Reset_h;
	 
	 
	 //Game state
	 GameState gamedata(.Clk, .Reset(Reset_h), .Frame_clk(VGA_VS), .Player_Attack(player_attack), .Player_X, .Player_Y, .Enemy1_X, .Enemy1_Y,
							  .Enemy2_X, .Enemy2_Y, .Enemy3_X, .Enemy3_Y, .Enemy4_X, .Enemy4_Y, .Enemy5_X, .Enemy5_Y,
							  .Damage_E1, .Damage_E2, .Damage_E3, .Damage_E4, .Damage_E5, 
								.health, .score1, .score2, .game_over);
	
	 EntityInterface entities(.select, .clk(Clk), .read, .write, .sel_dir,
										.Enemy1_X, .Enemy2_X, .Enemy3_X, .Enemy4_X, .Enemy5_X, .Player_X,
										.Enemy1_Y, .Enemy2_Y, .Enemy3_Y, .Enemy4_Y, .Enemy5_Y, .Player_Y,
										.Enemy1_Active, .Enemy2_Active, .Enemy3_Active, .Enemy4_Active, .Enemy5_Active,
										.Type_E1, .Type_E2, .Type_E3, .Type_E4, .Type_E5,
										.toNIOS_X, .toNIOS_Y, .toNIOS_Type,
										.toEnemy1_dir, .toEnemy2_dir, .toEnemy3_dir, .toEnemy4_dir, .toEnemy5_dir,
										.toNIOS_Active);
	 
	 //Level Data
	 level_rom level_instance(.DrawX, .DrawY, .room, .bg_type);
	 RoomState room_logic(.doorcode, .vsync(VGA_VS), .Reset(game_reset), .room, .initialize_room(initialize));
	 
	 //Draw modules
	 Background bg(.Red(bg_r), .Green(bg_g), .Blue(bg_b), 
						.bg_type, .DrawX, .DrawY);
						
	 TextDisplay text(.DrawX, .DrawY, .is_drawn(draw_text), .score1, .score2, .health,
							.addr(font_addr), .offset(text_offset));
							
	 Player player_instance(.Clk, .Reset(game_reset), .frame_clk(VGA_VS), .room, .doorcode,
									.keycode(keycode[7:0]), .Player_X, .Player_Y, .attack(player_attack));
	 
	 //Five enemies
	 Enemy enemy1(.Reset(game_reset), .frame_clk(VGA_VS), .Clk, .damage(Damage_E1), .initialize, .dir(toEnemy1_dir), .room, .number(3'b001),
						.Enemy_X(Enemy1_X), .Enemy_Y(Enemy1_Y), .active(Enemy1_Active), .Enemy_Type(Type_E1));
						
	 Enemy enemy2(.Reset(game_reset), .frame_clk(VGA_VS), .Clk, .damage(Damage_E2), .initialize, .dir(toEnemy2_dir), .room, .number(3'b010),
						.Enemy_X(Enemy2_X), .Enemy_Y(Enemy2_Y), .active(Enemy2_Active), .Enemy_Type(Type_E2));
						
	 Enemy enemy3(.Reset(game_reset), .frame_clk(VGA_VS), .Clk, .damage(Damage_E3), .initialize, .dir(toEnemy3_dir), .room, .number(3'b011),
						.Enemy_X(Enemy3_X), .Enemy_Y(Enemy3_Y), .active(Enemy3_Active), .Enemy_Type(Type_E3));
						
	 Enemy enemy4(.Reset(game_reset), .frame_clk(VGA_VS), .Clk, .damage(Damage_E4), .initialize, .dir(toEnemy4_dir), .room, .number(3'b100),
						.Enemy_X(Enemy4_X), .Enemy_Y(Enemy4_Y), .active(Enemy4_Active), .Enemy_Type(Type_E4));
						
	 Enemy enemy5(.Reset(game_reset), .frame_clk(VGA_VS), .Clk, .damage(Damage_E5), .initialize, .dir(toEnemy5_dir), .room, .number(3'b101),
						.Enemy_X(Enemy5_X), .Enemy_Y(Enemy5_Y), .active(Enemy5_Active), .Enemy_Type(Type_E5));
	 
	 //Interface modules
    VGA_controller vga_controller_instance(.Clk, 
														.Reset(Reset_h), 
														.VGA_HS, 
														.VGA_VS,
														.VGA_CLK,
														.VGA_BLANK_N,
														.VGA_SYNC_N,
														.DrawX,
														.DrawY);
    
    
    color_mapper color_instance(.DrawX,
										  .DrawY,
										  .Player_X, .Player_Y,
										  .Enemy1_X, .Enemy1_Y,
										  .Enemy2_X, .Enemy2_Y,
										  .Enemy3_X, .Enemy3_Y,
										  .Enemy4_X, .Enemy4_Y,
										  .Enemy5_X, .Enemy5_Y,
										  .E1_Type(Type_E1), .E2_Type(Type_E2), .E3_Type(Type_E3), .E4_Type(Type_E4), .E5_Type(Type_E5),
										  .frame_clk(VGA_VS), .player_attack,
										  .bg_r, .bg_g, .bg_b,
										  .font_addr, .text_offset, .draw_text,
										  .VGA_R,
										  .VGA_G,
										  .VGA_B);
    
    // Display keycode on hex display
    HexDriver hex_inst_0 (keycode[3:0], HEX0);
    HexDriver hex_inst_1 (keycode[7:4], HEX1);
    
endmodule
