module sprite_rom ( input [9:0]	addr,
						output [31:0]	data
					 );

	parameter SPRITE_NUMBER = 18;
   parameter DATA_WIDTH =  32;
				
	// ROM definition				
	parameter [0:32*SPRITE_NUMBER][DATA_WIDTH-1:0] ROM = {
		  //Wall Tile, code 0
        32'b11111111111111111111111111111111,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b11111111111111111111111111111111,
		  
		  //Floor Tile, code 1
		  32'b00000000000000000000000000000000,
		  32'b00000111111111111111111111100000,
		  32'b00011111111111111111111111111000,
		  32'b00100000000000000000000000000100,
		  32'b00101111111111111111111111110100,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b00101111111111111111111111110100,
		  32'b00100000000000000000000000000100,
		  32'b00011111111111111111111111111000,
		  32'b00000111111111111111111111100000,
		  32'b00000000000000000000000000000000,
		  
		  //BASE 2
		  //PLAYER OUTLINE 1
		   32'b00000000000011111111000000000000,
			32'b00000000000111111111100000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000000111111111100000000000,
			32'b00011100000011111111000000111000,
			32'b01111111100000111100000111111110,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111011111111111111111111011111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b01100011111111111111111111000110,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000001111111111111111110000000,
			32'b00000001111111111111111110000000,
			32'b00000001111111111111111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000000000000000000,
			
			
			//BASE 3
			//PLAYER COLOR 1
			32'b00000000000011111111000000000000,
			32'b00000000000111111111100000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000000111111111100000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000001111110000000000000,
			32'b00000000000000111100000000000000,
			32'b00011100000000011000000000111000,
			32'b01111111100000000000000111111110,
			32'b01111111111111000011111111111110,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111011111111111111111111011111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000001111111111111111110000000,
			32'b00000000011111111111111000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000000000000000000,
			
			
			//BASE 4
			//PLAYER OUTLINE 2
			32'b00000000000011111111000000000000,
			32'b00000000000111111111100000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000000111111111100000000000,
			32'b00011100000011111111000000111000,
			32'b01111111100000111100000111111110,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111011111111111111111111011111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b01100011111111111111111111000110,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000001111111111111111110000000,
			32'b00000001111111111111111110000000,
			32'b00000001111111111111111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000000000000000001111110000000,
			
			
			//BASE 5
			//PLAYER COLOR 2
			32'b00000000000011111111000000000000,
			32'b00000000000111111111100000000000,
			32'b00000000001111111111110000000000,
			32'b00000000001111111111110000000000,
			32'b00000000000111111111100000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000001111110000000000000,
			32'b00000000000000111100000000000000,
			32'b00011100000000011000000000111000,
			32'b01111111100000000000000111111110,
			32'b01111111111111000011111111111110,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111111111111111111111111111111,
			32'b11111011111111111111111111011111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000001111111111111111110000000,
			32'b00000000011111111111111000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000000000000000000000000,
			32'b00000001111110000000000000000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000000000000000001111110000000,
			
			
			//BASE 6
			//PLAYER OUTLINE ATTACK
			32'b00000000000011111111000111000000,
			32'b00000000000111111111100011101100,
			32'b00000000001111111111110001111100,
			32'b00000000001111111111110000111000,
			32'b00000000001111111111110001111100,
			32'b00000000001111111111110001101100,
			32'b00000000001111111111110000001100,
			32'b00000000000111111111100000011110,
			32'b00011100000011111111000000111110,
			32'b01111111100000111100000111111110,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111110,
			32'b11111111111111111111111111111110,
			32'b11111111111111111111111111111000,
			32'b11111111111111111111111111100000,
			32'b11111011111111111111111111000000,
			32'b11110011111111111111111111000000,
			32'b11110011111111111111111111000000,
			32'b11110011111111111111111111000000,
			32'b11110011111111111111111111000000,
			32'b01100011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000001111111111111111110000000,
			32'b00000001111111111111111110000000,
			32'b00000001111111111111111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000000000000000001111110000000,
			
			
			//BASE 7
			//PLAYER COLOR ATTACK
			32'b00000000000011111111000111000000,
			32'b00000000000111111111100011101100,
			32'b00000000001111111111110001111100,
			32'b00000000001111111111110000111000,
			32'b00000000000111111111100001111100,
			32'b00000000000011111111000001101100,
			32'b00000000000001111110000000000000,
			32'b00000000000000111100000000000000,
			32'b00011100000000011000000000111110,
			32'b01111111100000000000000111111110,
			32'b01111111111111000011111111111110,
			32'b11111111111111111111111111111110,
			32'b11111111111111111111111111111110,
			32'b11111111111111111111111111111000,
			32'b11111111111111111111111111100000,
			32'b11111011111111111111111111000000,
			32'b11110011111111111111111111000000,
			32'b11110011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000001111111111111111110000000,
			32'b00000000011111111111111000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000000000000000000000000,
			32'b00000001111110000000000000000000,
			32'b00000001111110000001111110000000,
			32'b00000001111110000001111110000000,
			32'b00000000000000000001111110000000,
			
			//BASE 8
			//KEESE OUTLINE 1
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b10000000000010000001000000000001,
			32'b11000000000011000011000000000011,
			32'b11100000000011100111000000000111,
			32'b11110000000011111111000000001111,
			32'b11111000000011111111000000011111,
			32'b01111000000011111111000000011110,
			32'b01111111000011111111000011111110,
			32'b01111111111011111111011111111110,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00011111111111111111111111111000,
			32'b00011111111111111111111111111000,
			32'b00011111111111111111111111111000,
			32'b00001111111111111111111111110000,
			32'b00001111111111111111111111110000,
			32'b00000111111111111111111111100000,
			32'b00000011111111111111111111000000,
			32'b00000000111111111111111100000000,
			32'b00000000000111111111100000000000,
			32'b00000000000001111110000000000000,
			32'b00000000000000111100000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			
			
			//BASE 9
			//KEESE COLOR 1
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b10000000000010000001000000000001,
			32'b11000000000011000011000000000011,
			32'b10100000000010100101000000000101,
			32'b10010000000010111101000000001001,
			32'b10001000000011000011000000010001,
			32'b01001000000010000001000000010010,
			32'b01000111000010100101000011100010,
			32'b01000000111010000001011100000010,
			32'b01000000000110000001100000000010,
			32'b00100000000010111101000000000100,
			32'b00100000000010100101000000000100,
			32'b00100000000010000001000000000100,
			32'b00100000000010000001000000000100,
			32'b00010000000010000001000000001000,
			32'b00010000000010000001000000001000,
			32'b00010000000010000001000000001000,
			32'b00001000000010000001000000010000,
			32'b00001000000010000001000000010000,
			32'b00000100000010000001000000100000,
			32'b00000011000010000001000011000000,
			32'b00000000111010000001011100000000,
			32'b00000000000110000001100000000000,
			32'b00000000000001000010000000000000,
			32'b00000000000000111100000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			
			
			//BASE 10
			//KEESE OUTLINE 2
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000010000001000000000000,
			32'b00000000000011000011000000000000,
			32'b00000000000011100111000000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000011111111000000000000,
			32'b00000000000111111111100000000000,
			32'b00000000111111111111111100000000,
			32'b00000011111111111111111111000000,
			32'b00000111111111111111111111100000,
			32'b00001111111111111111111111110000,
			32'b00001111111111111111111111110000,
			32'b00011111111111111111111111111000,
			32'b00011111111111111111111111111000,
			32'b00011111111111111111111111111000,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b01111111111001111110011111111110,
			32'b01111111000000111100000011111110,
			32'b01111000000000000000000000011110,
			32'b11111000000000000000000000011111,
			32'b11110000000000000000000000001111,
			32'b11100000000000000000000000000111,
			32'b11000000000000000000000000000011,
			32'b10000000000000000000000000000001,
			
			
			//BASE 11
			//KEESE COLOR 2
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000010000001000000000000,
			32'b00000000000011000011000000000000,
			32'b00000000000010100101000000000000,
			32'b00000000000010111101000000000000,
			32'b00000000000011000011000000000000,
			32'b00000000000010000001000000000000,
			32'b00000000000010100101000000000000,
			32'b00000000000010000001000000000000,
			32'b00000000000110000001100000000000,
			32'b00000000111010111101011100000000,
			32'b00000011000010100101000011000000,
			32'b00000100000010000001000000100000,
			32'b00001000000010000001000000010000,
			32'b00001000000010000001000000010000,
			32'b00010000000010000001000000001000,
			32'b00010000000010000001000000001000,
			32'b00010000000010000001000000001000,
			32'b00100000000010000001000000000100,
			32'b00100000000010000001000000000100,
			32'b00100000000010000001000000000100,
			32'b00100000000010000001000000000100,
			32'b01000000000110000001100000000010,
			32'b01000000111001000010011100000010,
			32'b01000111000000111100000011100010,
			32'b01001000000000000000000000010010,
			32'b10001000000000000000000000010001,
			32'b10010000000000000000000000001001,
			32'b10100000000000000000000000000101,
			32'b11000000000000000000000000000011,
			32'b10000000000000000000000000000001,
			
			//BASE 12
			//ZOMBIE OUTLINE 1
			32'b00000000000000000000000000000000,
			32'b00000000000001000000000000000000,
			32'b00000000000001101000000000000000,
			32'b00000000000001111100000000000000,
			32'b00000000011111111111111000000000,
			32'b00000011111111111111111111000000,
			32'b00000111111111111111111111100000,
			32'b00001111111111111111111111110000,
			32'b00011111111111111111111111111000,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b01111111111111111111111111111110,
			32'b11110111111111111111111111101111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b11110111111111111111111111101111,
			32'b00000111111111111111111111100000,
			32'b00000111111111111111111111100000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000111111111111111111111100000,
			32'b00000111111111111111111111100000,
			32'b00000111111111111111111111100000,
			32'b00001111111111111111111111110000,
			32'b00001111111111100111111111110000,
			32'b00001111111111000011111111110000,
			32'b00001111111110000001111111110000,
			32'b00001111110000000000001111110000,
			32'b00001111110000000000001111110000,
			32'b00001111110000000000000000000000,
			
			
			//BASE 13
			//ZOMBIE COLOR 1
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000011100000000111000000000,
			32'b00000011111111111111111111000000,
			32'b00000110111111111111100101100000,
			32'b00001100111111111111101100110000,
			32'b00011000111111111111100100011000,
			32'b00110001110111111111000110001100,
			32'b00100011100111111110011111000100,
			32'b00100111100111111110111111100100,
			32'b01000111101111111111111111100010,
			32'b01001111111111111111111111110010,
			32'b10010111111110111111111111101001,
			32'b10010011111110000011111001001001,
			32'b10010011111111111011110011001001,
			32'b11110111111111111111110111101111,
			32'b00000111111111111111100111100000,
			32'b00000110111111111111111101100000,
			32'b00000011000011100111000011000000,
			32'b00000011111100000000111111000000,
			32'b00000111111111111111111111100000,
			32'b00000111011111111111100011100000,
			32'b00000110011111111111110011100000,
			32'b00001110111111111111110000110000,
			32'b00001100111011100111111100110000,
			32'b00001111111011000011111110010000,
			32'b00001111111110000001111111110000,
			32'b00001000010000000000001000010000,
			32'b00001000010000000000001111110000,
			32'b00001111110000000000000000000000,
			
			
			//BASE 14
			//ZOMBIE OUTLINE 2
			32'b00000000000000000000000000000000,
			32'b00000000000001000000000000000000,
			32'b00000000000001101000000000000000,
			32'b00000000000001111100000000000000,
			32'b00000000011111111111111000000000,
			32'b00000011111111111111111111000000,
			32'b00000111111111111111111111100000,
			32'b00001111111111111111111111110000,
			32'b00011111111111111111111111111000,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b01111111111111111111111111111110,
			32'b11110111111111111111111111101111,
			32'b11110011111111111111111111001111,
			32'b11110011111111111111111111001111,
			32'b11110111111111111111111111101111,
			32'b00000111111111111111111111100000,
			32'b00000111111111111111111111100000,
			32'b00000011111111111111111111000000,
			32'b00000011111111111111111111000000,
			32'b00000111111111111111111111100000,
			32'b00000111111111111111111111100000,
			32'b00000111111111111111111111100000,
			32'b00001111111111111111111111110000,
			32'b00001111111111100111111111110000,
			32'b00001111111111000011111111110000,
			32'b00001111111110000001111111110000,
			32'b00001111110000000000001111110000,
			32'b00001111110000000000001111110000,
			32'b00000000000000000000001111110000,
			
			
			//BASE 15
			//ZOMBIE COLOR 2
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b00000000011100000000111000000000,
			32'b00000011111111111111111111000000,
			32'b00000110111111111111100101100000,
			32'b00001100111111111111101100110000,
			32'b00011000111111111111100100011000,
			32'b00110001110111111111000110001100,
			32'b00100011100111111110011111000100,
			32'b00100111100111111110111111100100,
			32'b01000111101111111111111111100010,
			32'b01001111111111111111111111110010,
			32'b10010111111110111111111111101001,
			32'b10010011111110000011111001001001,
			32'b10010011111111111011110011001001,
			32'b11110111111111111111110111101111,
			32'b00000111111111111111100111100000,
			32'b00000110111111111111111101100000,
			32'b00000011000011100111000011000000,
			32'b00000011111100000000111111000000,
			32'b00000111111111111111111111100000,
			32'b00000111011111111111100011100000,
			32'b00000110011111111111110011100000,
			32'b00001110111111111111110000110000,
			32'b00001100111011100111111100110000,
			32'b00001111111011000011111110010000,
			32'b00001111111110000001111111110000,
			32'b00001000010000000000001000010000,
			32'b00001111110000000000001000010000,
			32'b00000000000000000000001111110000,
		
	
			//BASE 16
			//SLIDER OUTLINE
			32'b00000100010001000010001000100000,
			32'b00001110111011100111011101110000,
			32'b00011111111111111111111111111000,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b01111111111111111111111111111110,
			32'b11111111111111111111111111111111,
			32'b01111111111111111111111111111110,
			32'b00111111111111111111111111111100,
			32'b00011111111111111111111111111000,
			32'b00001110111011100111011101110000,
			32'b00000100010001000010001000100000,
			
			
			//BASE 17
			//SLIDER COLOR
			32'b00000100010001000010001000100000,
			32'b00001010101010100101010101010000,
			32'b00010001000100011000100010001000,
			32'b00111111111111111111111111111100,
			32'b01011000000000000000000000011010,
			32'b10010111110000000000001111101001,
			32'b01010100000000000000000000101010,
			32'b00110100000000000000000000101100,
			32'b01010100000000000000000000101010,
			32'b10010100000000000000000000101001,
			32'b01010000000000000000000000001010,
			32'b00110000000000000000000000001100,
			32'b01010000000000000000000000001010,
			32'b10010000000000000000000000001001,
			32'b01010000000000000000000000001010,
			32'b00110000000000000000000000001100,
			32'b00110000000000000000000000001100,
			32'b01010000000000000000000000001010,
			32'b10010000000000000000000000001001,
			32'b01010000000000000000000000001010,
			32'b00110000000000000000000000001100,
			32'b01010000000000000000000000001010,
			32'b10010100000000000000000000101001,
			32'b01010100000000000000000000101010,
			32'b00110100000000000000000000101100,
			32'b01010100000000000000000000101010,
			32'b10010111110000000000001111101001,
			32'b01011000000000000000000000011010,
			32'b00111111111111111111111111111100,
			32'b00010001000100011000100010001000,
			32'b00001010101010100101010101010000,
			32'b00000100010001000010001000100000
        };

	assign data = ROM[addr];

endmodule  