/*
Modified sprite table ROM
takes the input of DrawX and DrawY and returns
if a floor or wall should be drawn
1 = draw wall
0 = draw floor
*/
module level_rom ( input [9:0]	DrawX, DrawY,
						 input logic [2:0] room,
						 output logic bg_type
					 );

	logic [19:0] data;
	
	// ROM definition		
	//Each room contains 20x15 background tiles
	parameter [0:29][19:0] ROM = {
	     //Room 0
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000100000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111,
		  
		  //Room 1
		  20'b00000000000000000000,
		  20'b11111111111111111111,
		  20'b10000000000000000001,
        20'b10000000000000000001,
		  20'b10000000100000000001,
		  20'b10000000100000000001,
		  20'b10000000100000000001,
		  20'b10001111111111000001,
		  20'b10000000100000000001,
		  20'b10000000100000000001,
		  20'b10000000100000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b10000000000000000001,
		  20'b11111111111111111111,
        };

	always_comb begin
		  
		data = ROM[15 * room + (DrawY/32)];
		bg_type = data[DrawX/32];
	
	end

endmodule