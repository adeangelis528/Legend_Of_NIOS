module sprite_rom ( input [5:0]	addr,
						output [31:0]	data
					 );

	parameter ADDR_WIDTH = 5;
   parameter DATA_WIDTH =  32;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  //Wall Tile
        32'b11111111111111111111111111111111,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b10000000000000000000000000000001,
		  32'b11111111111111111111111111111111,
		  
		  //Floor Tile
		  32'b00000000000000000000000000000000,
		  32'b00000111111110000001111111100000,
		  32'b00011111111111111111111111111000,
		  32'b00100000000000000000000000000100,
		  32'b00101111111111000011111111110100,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111100111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b00101111111111100111111111110100,
		  32'b00100111111111011011111111100100,
		  32'b00100110111110100101111101100100,
		  32'b00100110111110100101111101100100,
		  32'b00100111111111011011111111100100,
		  32'b00101111111111100111111111110100,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111100111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b01101111111111111111111111110110,
		  32'b00101111111111000011111111110100,
		  32'b00100000000000000000000000000100,
		  32'b00011111111111111111111111111000,
		  32'b00000111111110000001111111100000,
		  32'b00000000000000000000000000000000,
        };

	assign data = ROM[addr];

endmodule  